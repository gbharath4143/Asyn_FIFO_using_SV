`include "FIFO.sv"

`include "com_fifo.sv"
`include "int_fifo.sv"
`include "txn_fifo.sv"

`include "sbd_fifo.sv"
`include "cov_fifo.sv"
`include "mon_fifo.sv"

`include "wr_bfm_fifo.sv"
`include "rd_bfm_fifo.sv"

`include "wr_gen_fifo.sv"
`include "rd_gen_fifo.sv"

`include "wr_age_fifo.sv"
`include "rd_age_fifo.sv"

`include "env_fifo.sv"

`include "top_fifo.sv"