`include "com_fifo.sv"

`include "FIFO.sv"

`include "int_fifo.sv"

`include "wr_txn_fifo.sv"
`include "rd_txn_fifo.sv"

`include "sbd_fifo.sv"

`include "wr_cov_fifo.sv"
`include "rd_cov_fifo.sv"

`include "wr_mon_fifo.sv"
`include "rd_mon_fifo.sv"

`include "wr_bfm_fifo.sv"
`include "rd_bfm_fifo.sv"

`include "wr_gen_fifo.sv"
`include "rd_gen_fifo.sv"

`include "wr_age_fifo.sv"
`include "rd_age_fifo.sv"

`include "env_fifo.sv"

`include "top_fifo.sv"
