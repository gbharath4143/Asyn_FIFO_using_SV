class wr_cov_fifo;
  task run();
    $display("COV");
  endtask  
endclass
